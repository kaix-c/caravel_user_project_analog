magic
tech sky130A
magscale 1 2
timestamp 1727974750
<< locali >>
rect 730 540 1330 610
rect 730 380 1000 540
rect 1290 380 1330 540
rect 730 190 1330 380
rect 730 -400 830 190
rect 1230 -400 1330 190
rect 730 -440 1330 -400
rect 730 -630 1330 -590
rect 730 -1210 830 -630
rect 1230 -1210 1330 -630
rect 730 -1380 1330 -1210
rect 730 -1540 1000 -1380
rect 1290 -1540 1330 -1380
rect 730 -1610 1330 -1540
<< viali >>
rect 1000 380 1290 540
rect 1000 -1540 1290 -1380
<< metal1 >>
rect 750 540 1310 590
rect 750 380 1000 540
rect 1290 380 1310 540
rect 750 330 1310 380
rect 900 -210 950 330
rect 460 -490 660 -420
rect 1000 -490 1050 80
rect 460 -540 1050 -490
rect 460 -620 660 -540
rect 900 -1330 950 -810
rect 1000 -1080 1050 -540
rect 1110 -490 1160 0
rect 1400 -490 1600 -420
rect 1110 -540 1600 -490
rect 1110 -1010 1160 -540
rect 1400 -620 1600 -540
rect 750 -1380 1310 -1330
rect 750 -1540 1000 -1380
rect 1290 -1540 1310 -1380
rect 750 -1590 1310 -1540
use sky130_fd_pr__nfet_g5v0d10v5_7DHE2Q  XM1
timestamp 1727970069
transform 1 0 1028 0 1 -908
box -278 -358 278 358
use sky130_fd_pr__pfet_g5v0d10v5_6HUAKP  XM2
timestamp 1727970069
transform 1 0 1028 0 1 -103
box -308 -397 308 397
<< labels >>
flabel metal1 780 360 980 560 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 780 -1560 980 -1360 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 460 -620 660 -420 0 FreeSans 256 0 0 0 VIN
port 1 nsew
flabel metal1 1400 -620 1600 -420 0 FreeSans 256 0 0 0 VOUT
port 2 nsew
<< end >>
