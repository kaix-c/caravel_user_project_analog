* NGSPICE file created from inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_g5v0d10v5_7DHE2Q a_50_n100# a_n242_n322# a_n108_n100# a_n50_n188#
X0 a_50_n100# a_n50_n188# a_n108_n100# a_n242_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6HUAKP a_n50_n197# a_50_n100# w_n308_n397# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n308_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt inverter VDD VIN VOUT VSS
XXM1 VOUT VSS VSS VIN sky130_fd_pr__nfet_g5v0d10v5_7DHE2Q
XXM2 VIN VOUT VDD VDD sky130_fd_pr__pfet_g5v0d10v5_6HUAKP
.ends

