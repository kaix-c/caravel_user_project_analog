** sch_path: /home/kai/efabless/inverter2/xschem/inverter.sch
.subckt inverter VDD VIN VOUT VSS
*.PININFO VIN:I VOUT:O VDD:B VSS:B
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends
.end
