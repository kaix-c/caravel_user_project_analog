** sch_path: /home/kai/efabless/xschem/inverter_tb.sch
**.subckt inverter_tb
x1 VDD VIN VOUT GND inverter
V1 VIN GND pulse(0 1.8 1ns 1ns 1ns 5ns 10ns)
V2 VDD GND 2.5
**** begin user architecture code


.tran 0.01n 1u
.saveall

.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/kai/efabless/xschem/inverter.sym
** sch_path: /home/kai/efabless/xschem/inverter.sch
.subckt inverter VDD VIN VOUT VSS
*.ipin VIN
*.opin VOUT
*.iopin VDD
*.iopin VSS
XM1 VOUT VIN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 VOUT VIN VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
